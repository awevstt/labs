library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

package lab2_3_Kostenko_pack is
    subtype my_logic is std_logic;
    type my_vector is array (integer range<>) of my_logic;

end package lab2_3_Kostenko_pack;
