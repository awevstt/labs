library ieee;
use ieee.std_logic_1164.all;

package lab2_2_Kostenko_pack is
    subtype my_logic is std_logic;

end package lab2_2_Kostenko_pack;
